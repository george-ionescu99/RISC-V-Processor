`timescale 1ns / 1ps



//module ID_EX_reg(clk, reset,
//                 PC_ID, INSTRUCTION_ID, IMM_ID, REG_DATA1_ID, REG_DATA2_ID,
//                 FUNCT3_ID, FUNCT7_ID, OPCODE_ID, RD_ID, RS1_ID, RS2_ID,
//                 RegWrite_ID, MemToReg_ID, MemRead_ID, MemWrite_ID, ALUop_ID, Branch_ID);
                 
//output [31:0] PC_ID,          //adresa PC a instructiunii din etapa ID
//output [31:0] INSTRUCTION_ID, //instructiunea curenta in etapa ID
//output [31:0] IMM_ID,         //valoarea calculata
//                    output [31:0] REG_DATA1_ID,   //valoarea primului registru sursa citit
//                    output [31:0] REG_DATA2_ID,   //valoarea celui de-al doilea registru sursa citit
                    
//                    output [2:0] FUNCT3_ID,  //funct3 din codificarea instructiunii
//                    output [6:0] FUNCT7_ID,  //funct7 din codificarea instructiunii
//                    output [6:0] OPCODE_ID,     //opcode-ul instructiunii
//                    output [4:0] RD_ID,      //registru destinatie
//                    output [4:0] RS1_ID,     //registru sursa1
//                    output [4:0] RS2_ID,    //registru sursa2 
                    
                    
//                    //semnalele de control generate in ID
//                    output RegWrite_ID,  //semnal pentru scrierea in bancul de registri
//                    output MemtoReg_ID,  //semnal pentru scrierea din memorie in registru
//                    output MemRead_ID,   //semnal pentru citirea din memoria de date
//                    output MemWrite_ID,  //semnal pentru scrierea in memoria de date
//                    output [1:0] ALUop_ID, //codificarea operatiei efectuate de ALU 
//                    output ALUSrc_ID,      //semnal pentru alegerea operanzilor in ALU
//                    output Branch_ID);     //semnal pentru instructiuni de salt                 
                 
//endmodule
